library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

entity hier_MCU_SPI is
  port (
    MCU_PLL_SPI_CLK : in STD_LOGIC;
    MCU_PLL_SPI_SDIO : in STD_LOGIC;
    MCU_SP7_PMCU_SPI_AFE_PLL_CS2 : in STD_LOGIC;
    MCU_SP7_PMCU_SPI_AFE_PLL_CS2_2V5 : out STD_LOGIC;
    MCU_SP7_PMCU_SPI_DIG_PLL_CS1 : in STD_LOGIC;
    MCU_SP7_PMCU_SPI_DIG_PLL_CS1_2V5 : out STD_LOGIC;
    SP7_PLL4_SPI_SCK_2V5 : out STD_LOGIC;
    SP7_PLL_SPI_SDIO_o : out STD_LOGIC;
    clk_10mhz : in STD_LOGIC;
    rstn_10mhz : in STD_LOGIC
  );
end hier_MCU_SPI;

architecture STRUCTURE of hier_MCU_SPI is

  component MCU_PLL_SPI is
  port (
    clk_10mhz : in STD_LOGIC;
    rstn_10mhz : in STD_LOGIC;
    MCU_PLL_SPI_CLK : in STD_LOGIC;
    MCU_PLL_SPI_SDIO_i : in STD_LOGIC;
    MCU_PLL1_SPI_CS1 : in STD_LOGIC;
    MCU_PLL2_SPI_CS2 : in STD_LOGIC;
    MCU_PLL3_SPI_CS3 : in STD_LOGIC;
    MCU_PLL4_SPI_CS0 : in STD_LOGIC;
    SP7_PLL_SPI_SDIO_o : out STD_LOGIC;
    SP7_PLL_SPI_CLK : out STD_LOGIC;
    SP7_PLL4_SPI_CS : out STD_LOGIC;
    SP7_PLL1_SPI_CS1 : out STD_LOGIC;
    SP7_PLL2_SPI_CS2 : out STD_LOGIC;
    SP7_PLL3_SPI_CS3 : out STD_LOGIC;
    SP7_PLL4_SPI_SDI : out STD_LOGIC;
    SP7_PLL4_SPI_SDO : in STD_LOGIC
  );
  end component;
  
  signal MCU_PLL1_SPI_CS1 : STD_LOGIC;
  signal MCU_PLL4_SPI_CS0 : STD_LOGIC;
  signal MCU_PLL_SPI_0_SP7_PLL_SPI_SDIO_o : STD_LOGIC;
  signal MCU_PLL_SPI_SDIO_i : STD_LOGIC;
  signal SP7_PLL1_SPI_CS1 : STD_LOGIC;
  signal SP7_PLL4_SPI_CS : STD_LOGIC;
  signal SP7_PLL_SPI_CLK : STD_LOGIC;
  signal clk_wiz_0_clk_10 : STD_LOGIC;
  signal rstn : STD_LOGIC;
  signal xlconstant_0_dout : STD_LOGIC_VECTOR ( 0 to 0 ) := "1";
  signal NLW_MCU_PLL_SPI_0_SP7_PLL2_SPI_CS2_UNCONNECTED : STD_LOGIC;
  signal NLW_MCU_PLL_SPI_0_SP7_PLL3_SPI_CS3_UNCONNECTED : STD_LOGIC;
  signal NLW_MCU_PLL_SPI_0_SP7_PLL4_SPI_SDI_UNCONNECTED : STD_LOGIC;
  
begin

  MCU_PLL1_SPI_CS1 <= MCU_SP7_PMCU_SPI_AFE_PLL_CS2;
  MCU_PLL4_SPI_CS0 <= MCU_SP7_PMCU_SPI_DIG_PLL_CS1;
  MCU_PLL_SPI_SDIO_i <= MCU_PLL_SPI_SDIO;
  MCU_SP7_PMCU_SPI_AFE_PLL_CS2_2V5 <= SP7_PLL1_SPI_CS1;
  MCU_SP7_PMCU_SPI_DIG_PLL_CS1_2V5 <= SP7_PLL4_SPI_CS;
  SP7_PLL4_SPI_SCK_2V5 <= SP7_PLL_SPI_CLK;
  SP7_PLL_SPI_SDIO_o <= MCU_PLL_SPI_0_SP7_PLL_SPI_SDIO_o;
  clk_wiz_0_clk_10 <= clk_10mhz;
  rstn <= rstn_10mhz;
  
MCU_PLL_SPI_0: component MCU_PLL_SPI
     port map (
      MCU_PLL1_SPI_CS1 => MCU_PLL1_SPI_CS1,
      MCU_PLL2_SPI_CS2 => xlconstant_0_dout(0),
      MCU_PLL3_SPI_CS3 => xlconstant_0_dout(0),
      MCU_PLL4_SPI_CS0 => MCU_PLL4_SPI_CS0,
      MCU_PLL_SPI_CLK => MCU_PLL_SPI_CLK,
      MCU_PLL_SPI_SDIO_i => MCU_PLL_SPI_SDIO_i,
      SP7_PLL1_SPI_CS1 => SP7_PLL1_SPI_CS1,
      SP7_PLL2_SPI_CS2 => NLW_MCU_PLL_SPI_0_SP7_PLL2_SPI_CS2_UNCONNECTED,
      SP7_PLL3_SPI_CS3 => NLW_MCU_PLL_SPI_0_SP7_PLL3_SPI_CS3_UNCONNECTED,
      SP7_PLL4_SPI_CS => SP7_PLL4_SPI_CS,
      SP7_PLL4_SPI_SDI => NLW_MCU_PLL_SPI_0_SP7_PLL4_SPI_SDI_UNCONNECTED,
      SP7_PLL4_SPI_SDO => xlconstant_0_dout(0),
      SP7_PLL_SPI_CLK => SP7_PLL_SPI_CLK,
      SP7_PLL_SPI_SDIO_o => MCU_PLL_SPI_0_SP7_PLL_SPI_SDIO_o,
      clk_10mhz => clk_wiz_0_clk_10,
      rstn_10mhz => rstn
    );

end STRUCTURE;