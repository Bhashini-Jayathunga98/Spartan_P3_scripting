library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
entity sp7_cal3_wrapper is
  port (
    AFE_PLL_SP7_CLKSEL0 : out STD_LOGIC;
    AFE_PLL_SP7_LOCK_STAT : in STD_LOGIC;
    AFE_VCXO_SP7_122M88_CLK_LVDS_N : in STD_LOGIC;
    AFE_VCXO_SP7_122M88_CLK_LVDS_P : in STD_LOGIC;
    DIG_PLL_SP7_CLKSEL0 : out STD_LOGIC;
    DIG_PLL_SP7_LOCK_STAT : in STD_LOGIC;
    DMCU_DEV_SPI_SP7_CS : in STD_LOGIC;
    DMCU_FAN_CTRL : in STD_LOGIC;
    DMCU_LS_PORESET_CMD : in STD_LOGIC;
    DMCU_MAIN_CLK_EN : in STD_LOGIC;
    DMCU_PLL_RESETB : in STD_LOGIC;
    DMCU_RX_SP7_TX_UART_GPIO : out STD_LOGIC_VECTOR ( 0 to 0 );
    DMCU_SP7_AUXB_CONFIG_CMD : out STD_LOGIC_VECTOR ( 0 to 0 );
    DMCU_SP7_PMCU_SPI_AFE_PLL_CS2 : in STD_LOGIC;
    DMCU_SP7_PMCU_SPI_CLK : in STD_LOGIC;
    DMCU_SP7_PMCU_SPI_DIG_PLL_CS1 : in STD_LOGIC;
    DMCU_SP7_PMCU_SPI_MOSI : in STD_LOGIC;
    DMCU_SP7_ZU_SPI_MISO : out STD_LOGIC;
    DMCU_SP7_ZU_SPI_MOSI : in STD_LOGIC;
    DMCU_SP7_ZU_SPI_SCK : in STD_LOGIC;
    DMCU_SYSTEM_READY : in STD_LOGIC;
    DMCU_TX_SP7_RX_UART_GPIO : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_1 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_2 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_3 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_4 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_5 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_6 : in STD_LOGIC;
    GNSS_1PPS : in STD_LOGIC;
    GNSS_TP2 : in STD_LOGIC;
    GNSS_UART_RXD_SP7_TXD : out STD_LOGIC;
    GNSS_UART_TXD_SP7_RXD : in STD_LOGIC;
    J4124 : out STD_LOGIC_VECTOR ( 0 to 0 );
    J4142 : out STD_LOGIC_VECTOR ( 0 to 0 );
    KU_GNSS_1PPS : out STD_LOGIC;
    LOC_10M_OSC_SP7_ENABLE : out STD_LOGIC;
    LS_2V5_DDR_PG : in STD_LOGIC;
    LS_DDR4_TERM_PG : in STD_LOGIC;
    LS_GNSS_1PPS : out STD_LOGIC;
    LS_GNSS_TP2_GPIO : out STD_LOGIC;
    LS_PWRSEQ_RST_OUT_B_1V8 : in STD_LOGIC;
    LS_SP7_ASLEEP : in STD_LOGIC;
    LS_SP7_DMCU_RESET_STAT : out STD_LOGIC;
    LS_SP7_HRESET_B : in STD_LOGIC;
    LS_SP7_RESET_REQ_B : in STD_LOGIC;
    LS_SP7_SPI_CS1 : in STD_LOGIC;
    LS_SPI_CLK : in STD_LOGIC;
    LS_SPI_MISO : inout STD_LOGIC;
    LS_SPI_MOSI : in STD_LOGIC;
    LS_TA_PROG_SFP_PG : in STD_LOGIC;
    OCXO_CLK_BUF_ENB : out STD_LOGIC;
    OCXO_SP7_10M_DET_N : in STD_LOGIC;
    OCXO_SP7_10M_DET_P : in STD_LOGIC;
    SP7_10MHZ_LVDS_CLK_IN_N : in STD_LOGIC;
    SP7_10MHZ_LVDS_CLK_IN_P : in STD_LOGIC;
    SP7_10M_CLK_DAC_RESET : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_DAC_SCLK : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_DAC_SDIN : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_DAC_SEL : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_DAC_SYNC : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_REF_EN_B : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_SOURCE_SEL : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_12V_OCXO_EN : out STD_LOGIC;
    SP7_3V3_AFEPLL_PG : in STD_LOGIC;
    SP7_3V3_DIGPLL_PG : in STD_LOGIC;
    SP7_3V3_OCXO_PG : in STD_LOGIC;
    SP7_3V3_VCXO_PG : in STD_LOGIC;
    SP7_50MHZ_OSC_INPUT : in STD_LOGIC;
    SP7_AFE_PLL_RESETB : out STD_LOGIC;
    SP7_AFE_PLL_SPI_CS1 : out STD_LOGIC;
    SP7_AFE_PLL_SYNC : out STD_LOGIC;
    SP7_AFE_VCXO_ENB : out STD_LOGIC;
    SP7_AUXB_CONFIG_CMD : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_AUXB_CONFIG_STAT : in STD_LOGIC;
    SP7_AUXB_PWR_EN : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_AUXB_PWR_STAT : in STD_LOGIC;
    SP7_AUXETH_PLL_GPIO1_OE : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_AUXETH_PLL_GPIO4_LOCK : in STD_LOGIC;
    SP7_AUXETH_PLL_HW_SW_CTRL : inout STD_LOGIC;
    SP7_AUXETH_PLL_RESET : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_DBG_UART_RX : in STD_LOGIC;
    SP7_DBG_UART_TX : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_DIG_PLL_RESET : out STD_LOGIC;
    SP7_DIG_PLL_SPI_CS0 : out STD_LOGIC;
    SP7_DIG_PLL_SYNC : out STD_LOGIC;
    SP7_DIP_SW_11 : in STD_LOGIC;
    SP7_DIP_SW_12 : in STD_LOGIC;
    SP7_DIP_SW_21 : in STD_LOGIC;
    SP7_DIP_SW_22 : in STD_LOGIC;
    SP7_DIP_SW_32 : in STD_LOGIC;
    SP7_DMCU_AUXB_CONFIG_STAT : in STD_LOGIC;
    SP7_DMCU_IRQ : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_FAN_PWM_CTRL_1 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_2 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_3 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_4 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_5 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_6 : out STD_LOGIC;
    SP7_FAN_PWR_CTRL_EN : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_GNSS_KU_UART_RX : out STD_LOGIC;
    SP7_GNSS_LS_UART_RX : in STD_LOGIC;
    SP7_GNSS_LS_UART_TX : out STD_LOGIC;
    SP7_GNSS_RST_B : out STD_LOGIC;
    SP7_GNSS_ZU_UART_RX : out STD_LOGIC;
    SP7_JTAG_BUF_EN : in STD_LOGIC;
    SP7_KU_QSPI_CFG_MAP : out STD_LOGIC;
    SP7_KU_SPARE1N_CLKN_LVDS : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_KU_SPARE1P_CLKP_LVDS : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_LS_BST_EN_2V5 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_LS_DDR_RESET_B : out STD_LOGIC;
    SP7_LS_EMMC_RESET_B : out STD_LOGIC;
    SP7_LS_IRQ : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_LS_NOR_PORESET : out STD_LOGIC;
    SP7_LS_PORESET_CMD_2V5 : out STD_LOGIC;
    SP7_LS_QSPI_CFG_MAP_2V5 : out STD_LOGIC;
    SP7_LS_TA_PROG_SFP_EN_2V5 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_MAIN_CLK_STAT : out STD_LOGIC;
    SP7_OCXO_INTB_EXT_REF : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_OSC_PWR_EN : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_PLL_PWR_EN : out STD_LOGIC;
    SP7_PLL_SPI_CLK : out STD_LOGIC;
    SP7_PLL_SPI_SDIO : out STD_LOGIC;
    SP7_PLL_STATUS : out STD_LOGIC;
    SP7_PUDC : in STD_LOGIC;
    SP7_SPARE_LED_2 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_SPARE_LED_3 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_SPARE_LED_4 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_3V3_GPIO_1 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_3V3_GPIO_2 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_3V3_GPIO_3 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_3V3_GPIO_5 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_MODE_SPARE_LED_1 : out STD_LOGIC;
    SP7_ZU_QSPI_CFG_MAP_2V5 : out STD_LOGIC;
    SP7_ZU_SPARE1N_CLKN_LVDS : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_SPARE1P_CLKP_LVDS : out STD_LOGIC_VECTOR ( 0 to 0 );
    ZU_BOOT_STATUS_2V5 : in STD_LOGIC;
    ZU_DONE_2V5 : in STD_LOGIC;
    ZU_ERROR_OUT_2V5 : in STD_LOGIC;
    ZU_ERROR_STATUS_2V5 : in STD_LOGIC;
    ZU_GNSS_1PPS : out STD_LOGIC;
    ZU_SP7_DMCU_RESET_STAT : out STD_LOGIC;
    spi_rtl_0_io0_io : inout STD_LOGIC;
    spi_rtl_0_io1_io : inout STD_LOGIC;
    spi_rtl_0_io2_io : inout STD_LOGIC;
    spi_rtl_0_io3_io : inout STD_LOGIC;
    spi_rtl_0_ss_io : inout STD_LOGIC_VECTOR ( 0 to 0 )
  );
end sp7_cal3_wrapper;

architecture STRUCTURE of sp7_cal3_wrapper is
  component sp7_cal3 is
  port (
    GNSS_UART_TXD_SP7_RXD : in STD_LOGIC;
    SP7_DIP_SW_11 : in STD_LOGIC;
    SP7_DIP_SW_12 : in STD_LOGIC;
    SP7_DIP_SW_21 : in STD_LOGIC;
    SP7_DIP_SW_22 : in STD_LOGIC;
    SP7_DIP_SW_32 : in STD_LOGIC;
    DIG_PLL_SP7_LOCK_STAT : in STD_LOGIC;
    AFE_PLL_SP7_LOCK_STAT : in STD_LOGIC;
    SP7_AUXB_PWR_STAT : in STD_LOGIC;
    SP7_AUXB_CONFIG_STAT : in STD_LOGIC;
    LS_DDR4_TERM_PG : in STD_LOGIC;
    LS_2V5_DDR_PG : in STD_LOGIC;
    LS_TA_PROG_SFP_PG : in STD_LOGIC;
    GNSS_1PPS : in STD_LOGIC;
    GNSS_TP2 : in STD_LOGIC;
    ZU_DONE_2V5 : in STD_LOGIC;
    ZU_ERROR_OUT_2V5 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_1 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_2 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_3 : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_4 : in STD_LOGIC;
    ZU_BOOT_STATUS_2V5 : in STD_LOGIC;
    ZU_ERROR_STATUS_2V5 : in STD_LOGIC;
    SP7_3V3_DIGPLL_PG : in STD_LOGIC;
    SP7_3V3_AFEPLL_PG : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_5 : in STD_LOGIC;
    SP7_3V3_OCXO_PG : in STD_LOGIC;
    SP7_3V3_VCXO_PG : in STD_LOGIC;
    FAN_SP7_TACH_SENSOR_6 : in STD_LOGIC;
    OCXO_SP7_10M_DET_P : in STD_LOGIC;
    OCXO_SP7_10M_DET_N : in STD_LOGIC;
    DMCU_MAIN_CLK_EN : in STD_LOGIC;
    DMCU_PLL_RESETB : in STD_LOGIC;
    LS_SP7_HRESET_B : in STD_LOGIC;
    LS_SP7_RESET_REQ_B : in STD_LOGIC;
    LS_SP7_ASLEEP : in STD_LOGIC;
    LS_SPI_MOSI : in STD_LOGIC;
    LS_SPI_CLK : in STD_LOGIC;
    LS_SP7_SPI_CS1 : in STD_LOGIC;
    DMCU_SP7_PMCU_SPI_MOSI : in STD_LOGIC;
    DMCU_SP7_PMCU_SPI_CLK : in STD_LOGIC;
    SP7_PUDC : in STD_LOGIC;
    DMCU_SYSTEM_READY : in STD_LOGIC;
    DMCU_SP7_ZU_SPI_SCK : in STD_LOGIC;
    DMCU_DEV_SPI_SP7_CS : in STD_LOGIC;
    DMCU_SP7_ZU_SPI_MOSI : in STD_LOGIC;
    SP7_GNSS_LS_UART_RX : in STD_LOGIC;
    SP7_DBG_UART_RX : in STD_LOGIC;
    LS_PWRSEQ_RST_OUT_B_1V8 : in STD_LOGIC;
    DMCU_LS_PORESET_CMD : in STD_LOGIC;
    DMCU_TX_SP7_RX_UART_GPIO : in STD_LOGIC;
    DMCU_FAN_CTRL : in STD_LOGIC;
    SP7_50MHZ_OSC_INPUT : in STD_LOGIC;
    DMCU_SP7_PMCU_SPI_AFE_PLL_CS2 : in STD_LOGIC;
    DMCU_SP7_PMCU_SPI_DIG_PLL_CS1 : in STD_LOGIC;
    SP7_GNSS_RST_B : out STD_LOGIC;
    GNSS_UART_RXD_SP7_TXD : out STD_LOGIC;
    SP7_SPARE_LED_2 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_SPARE_LED_3 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_SPARE_LED_4 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_REF_EN_B : out STD_LOGIC_VECTOR ( 0 to 0 );
    OCXO_CLK_BUF_ENB : out STD_LOGIC;
    SP7_10M_CLK_DAC_SEL : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_DAC_RESET : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_DAC_SDIN : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_DAC_SCLK : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_CLK_DAC_SYNC : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_DIG_PLL_SPI_CS0 : out STD_LOGIC;
    SP7_AFE_PLL_SPI_CS1 : out STD_LOGIC;
    SP7_PLL_SPI_CLK : out STD_LOGIC;
    SP7_KU_QSPI_CFG_MAP : out STD_LOGIC;
    SP7_AUXB_PWR_EN : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_AFE_VCXO_ENB : out STD_LOGIC;
    SP7_OSC_PWR_EN : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_DMCU_IRQ : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_MAIN_CLK_STAT : out STD_LOGIC;
    SP7_ZU_SPARE1P_CLKP_LVDS : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_KU_SPARE1P_CLKP_LVDS : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_DIG_PLL_SYNC : out STD_LOGIC;
    SP7_AFE_PLL_RESETB : out STD_LOGIC;
    SP7_AFE_PLL_SYNC : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_5 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_4 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_6 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_1 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_2 : out STD_LOGIC;
    SP7_FAN_PWM_CTRL_3 : out STD_LOGIC;
    SP7_DIG_PLL_RESET : out STD_LOGIC;
    SP7_LS_BST_EN_2V5 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_QSPI_CFG_MAP_2V5 : out STD_LOGIC;
    SP7_LS_QSPI_CFG_MAP_2V5 : out STD_LOGIC;
    SP7_FAN_PWR_CTRL_EN : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_LS_TA_PROG_SFP_EN_2V5 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_12V_OCXO_EN : out STD_LOGIC;
    SP7_LS_PORESET_CMD_2V5 : out STD_LOGIC;
    SP7_ZU_SPARE1N_CLKN_LVDS : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_KU_SPARE1N_CLKN_LVDS : out STD_LOGIC_VECTOR ( 0 to 0 );
    LS_SP7_DMCU_RESET_STAT : out STD_LOGIC;
    SP7_OCXO_INTB_EXT_REF : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_LS_IRQ : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_PLL_STATUS : out STD_LOGIC;
    SP7_LS_NOR_PORESET : out STD_LOGIC;
    SP7_LS_DDR_RESET_B : out STD_LOGIC;
    SP7_LS_EMMC_RESET_B : out STD_LOGIC;
    DMCU_SP7_ZU_SPI_MISO : out STD_LOGIC;
    ZU_SP7_DMCU_RESET_STAT : out STD_LOGIC;
    SP7_GNSS_LS_UART_TX : out STD_LOGIC;
    SP7_GNSS_KU_UART_RX : out STD_LOGIC;
    SP7_GNSS_ZU_UART_RX : out STD_LOGIC;
    SP7_ZU_MODE_SPARE_LED_1 : out STD_LOGIC;
    SP7_DBG_UART_TX : out STD_LOGIC_VECTOR ( 0 to 0 );
    DMCU_RX_SP7_TX_UART_GPIO : out STD_LOGIC_VECTOR ( 0 to 0 );
    LS_GNSS_1PPS : out STD_LOGIC;
    LS_GNSS_TP2_GPIO : out STD_LOGIC;
    KU_GNSS_1PPS : out STD_LOGIC;
    ZU_GNSS_1PPS : out STD_LOGIC;
    SP7_AUXB_CONFIG_CMD : out STD_LOGIC_VECTOR ( 0 to 0 );
    AFE_PLL_SP7_CLKSEL0 : out STD_LOGIC;
    DIG_PLL_SP7_CLKSEL0 : out STD_LOGIC;
    SP7_PLL_SPI_SDIO : out STD_LOGIC;
    SP7_DMCU_AUXB_CONFIG_STAT : in STD_LOGIC;
    DMCU_SP7_AUXB_CONFIG_CMD : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_AUXETH_PLL_RESET : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_AUXETH_PLL_GPIO4_LOCK : in STD_LOGIC;
    SP7_AUXETH_PLL_GPIO1_OE : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_10M_SOURCE_SEL : out STD_LOGIC_VECTOR ( 0 to 0 );
    LS_SPI_MISO : inout STD_LOGIC;
    J4124 : out STD_LOGIC_VECTOR ( 0 to 0 );
    J4142 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_3V3_GPIO_1 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_3V3_GPIO_5 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_3V3_GPIO_2 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_ZU_3V3_GPIO_3 : out STD_LOGIC_VECTOR ( 0 to 0 );
    SP7_JTAG_BUF_EN : in STD_LOGIC;
    SP7_10MHZ_LVDS_CLK_IN_P : in STD_LOGIC;
    SP7_10MHZ_LVDS_CLK_IN_N : in STD_LOGIC;
    AFE_VCXO_SP7_122M88_CLK_LVDS_P : in STD_LOGIC;
    AFE_VCXO_SP7_122M88_CLK_LVDS_N : in STD_LOGIC;
    LOC_10M_OSC_SP7_ENABLE : out STD_LOGIC;
    SP7_PLL_PWR_EN : out STD_LOGIC;
    SP7_AUXETH_PLL_HW_SW_CTRL : inout STD_LOGIC;
    spi_rtl_0_io0_i : in STD_LOGIC;
    spi_rtl_0_io0_o : out STD_LOGIC;
    spi_rtl_0_io0_t : out STD_LOGIC;
    spi_rtl_0_io1_i : in STD_LOGIC;
    spi_rtl_0_io1_o : out STD_LOGIC;
    spi_rtl_0_io1_t : out STD_LOGIC;
    spi_rtl_0_io2_i : in STD_LOGIC;
    spi_rtl_0_io2_o : out STD_LOGIC;
    spi_rtl_0_io2_t : out STD_LOGIC;
    spi_rtl_0_io3_i : in STD_LOGIC;
    spi_rtl_0_io3_o : out STD_LOGIC;
    spi_rtl_0_io3_t : out STD_LOGIC;
    spi_rtl_0_ss_i : in STD_LOGIC_VECTOR ( 0 to 0 );
    spi_rtl_0_ss_o : out STD_LOGIC_VECTOR ( 0 to 0 );
    spi_rtl_0_ss_t : out STD_LOGIC
  );
  end component sp7_cal3;
  component IOBUF is
  port (
    I : in STD_LOGIC;
    O : out STD_LOGIC;
    T : in STD_LOGIC;
    IO : inout STD_LOGIC
  );
  end component IOBUF;
  signal spi_rtl_0_io0_i : STD_LOGIC;
  signal spi_rtl_0_io0_o : STD_LOGIC;
  signal spi_rtl_0_io0_t : STD_LOGIC;
  signal spi_rtl_0_io1_i : STD_LOGIC;
  signal spi_rtl_0_io1_o : STD_LOGIC;
  signal spi_rtl_0_io1_t : STD_LOGIC;
  signal spi_rtl_0_io2_i : STD_LOGIC;
  signal spi_rtl_0_io2_o : STD_LOGIC;
  signal spi_rtl_0_io2_t : STD_LOGIC;
  signal spi_rtl_0_io3_i : STD_LOGIC;
  signal spi_rtl_0_io3_o : STD_LOGIC;
  signal spi_rtl_0_io3_t : STD_LOGIC;
  signal spi_rtl_0_ss_i_0 : STD_LOGIC_VECTOR ( 0 to 0 );
  signal spi_rtl_0_ss_io_0 : STD_LOGIC_VECTOR ( 0 to 0 );
  signal spi_rtl_0_ss_o_0 : STD_LOGIC_VECTOR ( 0 to 0 );
  signal spi_rtl_0_ss_t : STD_LOGIC;
begin
sp7_cal3_i: component sp7_cal3
     port map (
      AFE_PLL_SP7_CLKSEL0 => AFE_PLL_SP7_CLKSEL0,
      AFE_PLL_SP7_LOCK_STAT => AFE_PLL_SP7_LOCK_STAT,
      AFE_VCXO_SP7_122M88_CLK_LVDS_N => AFE_VCXO_SP7_122M88_CLK_LVDS_N,
      AFE_VCXO_SP7_122M88_CLK_LVDS_P => AFE_VCXO_SP7_122M88_CLK_LVDS_P,
      DIG_PLL_SP7_CLKSEL0 => DIG_PLL_SP7_CLKSEL0,
      DIG_PLL_SP7_LOCK_STAT => DIG_PLL_SP7_LOCK_STAT,
      DMCU_DEV_SPI_SP7_CS => DMCU_DEV_SPI_SP7_CS,
      DMCU_FAN_CTRL => DMCU_FAN_CTRL,
      DMCU_LS_PORESET_CMD => DMCU_LS_PORESET_CMD,
      DMCU_MAIN_CLK_EN => DMCU_MAIN_CLK_EN,
      DMCU_PLL_RESETB => DMCU_PLL_RESETB,
      DMCU_RX_SP7_TX_UART_GPIO(0) => DMCU_RX_SP7_TX_UART_GPIO(0),
      DMCU_SP7_AUXB_CONFIG_CMD(0) => DMCU_SP7_AUXB_CONFIG_CMD(0),
      DMCU_SP7_PMCU_SPI_AFE_PLL_CS2 => DMCU_SP7_PMCU_SPI_AFE_PLL_CS2,
      DMCU_SP7_PMCU_SPI_CLK => DMCU_SP7_PMCU_SPI_CLK,
      DMCU_SP7_PMCU_SPI_DIG_PLL_CS1 => DMCU_SP7_PMCU_SPI_DIG_PLL_CS1,
      DMCU_SP7_PMCU_SPI_MOSI => DMCU_SP7_PMCU_SPI_MOSI,
      DMCU_SP7_ZU_SPI_MISO => DMCU_SP7_ZU_SPI_MISO,
      DMCU_SP7_ZU_SPI_MOSI => DMCU_SP7_ZU_SPI_MOSI,
      DMCU_SP7_ZU_SPI_SCK => DMCU_SP7_ZU_SPI_SCK,
      DMCU_SYSTEM_READY => DMCU_SYSTEM_READY,
      DMCU_TX_SP7_RX_UART_GPIO => DMCU_TX_SP7_RX_UART_GPIO,
      FAN_SP7_TACH_SENSOR_1 => FAN_SP7_TACH_SENSOR_1,
      FAN_SP7_TACH_SENSOR_2 => FAN_SP7_TACH_SENSOR_2,
      FAN_SP7_TACH_SENSOR_3 => FAN_SP7_TACH_SENSOR_3,
      FAN_SP7_TACH_SENSOR_4 => FAN_SP7_TACH_SENSOR_4,
      FAN_SP7_TACH_SENSOR_5 => FAN_SP7_TACH_SENSOR_5,
      FAN_SP7_TACH_SENSOR_6 => FAN_SP7_TACH_SENSOR_6,
      GNSS_1PPS => GNSS_1PPS,
      GNSS_TP2 => GNSS_TP2,
      GNSS_UART_RXD_SP7_TXD => GNSS_UART_RXD_SP7_TXD,
      GNSS_UART_TXD_SP7_RXD => GNSS_UART_TXD_SP7_RXD,
      J4124(0) => J4124(0),
      J4142(0) => J4142(0),
      KU_GNSS_1PPS => KU_GNSS_1PPS,
      LOC_10M_OSC_SP7_ENABLE => LOC_10M_OSC_SP7_ENABLE,
      LS_2V5_DDR_PG => LS_2V5_DDR_PG,
      LS_DDR4_TERM_PG => LS_DDR4_TERM_PG,
      LS_GNSS_1PPS => LS_GNSS_1PPS,
      LS_GNSS_TP2_GPIO => LS_GNSS_TP2_GPIO,
      LS_PWRSEQ_RST_OUT_B_1V8 => LS_PWRSEQ_RST_OUT_B_1V8,
      LS_SP7_ASLEEP => LS_SP7_ASLEEP,
      LS_SP7_DMCU_RESET_STAT => LS_SP7_DMCU_RESET_STAT,
      LS_SP7_HRESET_B => LS_SP7_HRESET_B,
      LS_SP7_RESET_REQ_B => LS_SP7_RESET_REQ_B,
      LS_SP7_SPI_CS1 => LS_SP7_SPI_CS1,
      LS_SPI_CLK => LS_SPI_CLK,
      LS_SPI_MISO => LS_SPI_MISO,
      LS_SPI_MOSI => LS_SPI_MOSI,
      LS_TA_PROG_SFP_PG => LS_TA_PROG_SFP_PG,
      OCXO_CLK_BUF_ENB => OCXO_CLK_BUF_ENB,
      OCXO_SP7_10M_DET_N => OCXO_SP7_10M_DET_N,
      OCXO_SP7_10M_DET_P => OCXO_SP7_10M_DET_P,
      SP7_10MHZ_LVDS_CLK_IN_N => SP7_10MHZ_LVDS_CLK_IN_N,
      SP7_10MHZ_LVDS_CLK_IN_P => SP7_10MHZ_LVDS_CLK_IN_P,
      SP7_10M_CLK_DAC_RESET(0) => SP7_10M_CLK_DAC_RESET(0),
      SP7_10M_CLK_DAC_SCLK(0) => SP7_10M_CLK_DAC_SCLK(0),
      SP7_10M_CLK_DAC_SDIN(0) => SP7_10M_CLK_DAC_SDIN(0),
      SP7_10M_CLK_DAC_SEL(0) => SP7_10M_CLK_DAC_SEL(0),
      SP7_10M_CLK_DAC_SYNC(0) => SP7_10M_CLK_DAC_SYNC(0),
      SP7_10M_CLK_REF_EN_B(0) => SP7_10M_CLK_REF_EN_B(0),
      SP7_10M_SOURCE_SEL(0) => SP7_10M_SOURCE_SEL(0),
      SP7_12V_OCXO_EN => SP7_12V_OCXO_EN,
      SP7_3V3_AFEPLL_PG => SP7_3V3_AFEPLL_PG,
      SP7_3V3_DIGPLL_PG => SP7_3V3_DIGPLL_PG,
      SP7_3V3_OCXO_PG => SP7_3V3_OCXO_PG,
      SP7_3V3_VCXO_PG => SP7_3V3_VCXO_PG,
      SP7_50MHZ_OSC_INPUT => SP7_50MHZ_OSC_INPUT,
      SP7_AFE_PLL_RESETB => SP7_AFE_PLL_RESETB,
      SP7_AFE_PLL_SPI_CS1 => SP7_AFE_PLL_SPI_CS1,
      SP7_AFE_PLL_SYNC => SP7_AFE_PLL_SYNC,
      SP7_AFE_VCXO_ENB => SP7_AFE_VCXO_ENB,
      SP7_AUXB_CONFIG_CMD(0) => SP7_AUXB_CONFIG_CMD(0),
      SP7_AUXB_CONFIG_STAT => SP7_AUXB_CONFIG_STAT,
      SP7_AUXB_PWR_EN(0) => SP7_AUXB_PWR_EN(0),
      SP7_AUXB_PWR_STAT => SP7_AUXB_PWR_STAT,
      SP7_AUXETH_PLL_GPIO1_OE(0) => SP7_AUXETH_PLL_GPIO1_OE(0),
      SP7_AUXETH_PLL_GPIO4_LOCK => SP7_AUXETH_PLL_GPIO4_LOCK,
      SP7_AUXETH_PLL_HW_SW_CTRL => SP7_AUXETH_PLL_HW_SW_CTRL,
      SP7_AUXETH_PLL_RESET(0) => SP7_AUXETH_PLL_RESET(0),
      SP7_DBG_UART_RX => SP7_DBG_UART_RX,
      SP7_DBG_UART_TX(0) => SP7_DBG_UART_TX(0),
      SP7_DIG_PLL_RESET => SP7_DIG_PLL_RESET,
      SP7_DIG_PLL_SPI_CS0 => SP7_DIG_PLL_SPI_CS0,
      SP7_DIG_PLL_SYNC => SP7_DIG_PLL_SYNC,
      SP7_DIP_SW_11 => SP7_DIP_SW_11,
      SP7_DIP_SW_12 => SP7_DIP_SW_12,
      SP7_DIP_SW_21 => SP7_DIP_SW_21,
      SP7_DIP_SW_22 => SP7_DIP_SW_22,
      SP7_DIP_SW_32 => SP7_DIP_SW_32,
      SP7_DMCU_AUXB_CONFIG_STAT => SP7_DMCU_AUXB_CONFIG_STAT,
      SP7_DMCU_IRQ(0) => SP7_DMCU_IRQ(0),
      SP7_FAN_PWM_CTRL_1 => SP7_FAN_PWM_CTRL_1,
      SP7_FAN_PWM_CTRL_2 => SP7_FAN_PWM_CTRL_2,
      SP7_FAN_PWM_CTRL_3 => SP7_FAN_PWM_CTRL_3,
      SP7_FAN_PWM_CTRL_4 => SP7_FAN_PWM_CTRL_4,
      SP7_FAN_PWM_CTRL_5 => SP7_FAN_PWM_CTRL_5,
      SP7_FAN_PWM_CTRL_6 => SP7_FAN_PWM_CTRL_6,
      SP7_FAN_PWR_CTRL_EN(0) => SP7_FAN_PWR_CTRL_EN(0),
      SP7_GNSS_KU_UART_RX => SP7_GNSS_KU_UART_RX,
      SP7_GNSS_LS_UART_RX => SP7_GNSS_LS_UART_RX,
      SP7_GNSS_LS_UART_TX => SP7_GNSS_LS_UART_TX,
      SP7_GNSS_RST_B => SP7_GNSS_RST_B,
      SP7_GNSS_ZU_UART_RX => SP7_GNSS_ZU_UART_RX,
      SP7_JTAG_BUF_EN => SP7_JTAG_BUF_EN,
      SP7_KU_QSPI_CFG_MAP => SP7_KU_QSPI_CFG_MAP,
      SP7_KU_SPARE1N_CLKN_LVDS(0) => SP7_KU_SPARE1N_CLKN_LVDS(0),
      SP7_KU_SPARE1P_CLKP_LVDS(0) => SP7_KU_SPARE1P_CLKP_LVDS(0),
      SP7_LS_BST_EN_2V5(0) => SP7_LS_BST_EN_2V5(0),
      SP7_LS_DDR_RESET_B => SP7_LS_DDR_RESET_B,
      SP7_LS_EMMC_RESET_B => SP7_LS_EMMC_RESET_B,
      SP7_LS_IRQ(0) => SP7_LS_IRQ(0),
      SP7_LS_NOR_PORESET => SP7_LS_NOR_PORESET,
      SP7_LS_PORESET_CMD_2V5 => SP7_LS_PORESET_CMD_2V5,
      SP7_LS_QSPI_CFG_MAP_2V5 => SP7_LS_QSPI_CFG_MAP_2V5,
      SP7_LS_TA_PROG_SFP_EN_2V5(0) => SP7_LS_TA_PROG_SFP_EN_2V5(0),
      SP7_MAIN_CLK_STAT => SP7_MAIN_CLK_STAT,
      SP7_OCXO_INTB_EXT_REF(0) => SP7_OCXO_INTB_EXT_REF(0),
      SP7_OSC_PWR_EN(0) => SP7_OSC_PWR_EN(0),
      SP7_PLL_PWR_EN => SP7_PLL_PWR_EN,
      SP7_PLL_SPI_CLK => SP7_PLL_SPI_CLK,
      SP7_PLL_SPI_SDIO => SP7_PLL_SPI_SDIO,
      SP7_PLL_STATUS => SP7_PLL_STATUS,
      SP7_PUDC => SP7_PUDC,
      SP7_SPARE_LED_2(0) => SP7_SPARE_LED_2(0),
      SP7_SPARE_LED_3(0) => SP7_SPARE_LED_3(0),
      SP7_SPARE_LED_4(0) => SP7_SPARE_LED_4(0),
      SP7_ZU_3V3_GPIO_1(0) => SP7_ZU_3V3_GPIO_1(0),
      SP7_ZU_3V3_GPIO_2(0) => SP7_ZU_3V3_GPIO_2(0),
      SP7_ZU_3V3_GPIO_3(0) => SP7_ZU_3V3_GPIO_3(0),
      SP7_ZU_3V3_GPIO_5(0) => SP7_ZU_3V3_GPIO_5(0),
      SP7_ZU_MODE_SPARE_LED_1 => SP7_ZU_MODE_SPARE_LED_1,
      SP7_ZU_QSPI_CFG_MAP_2V5 => SP7_ZU_QSPI_CFG_MAP_2V5,
      SP7_ZU_SPARE1N_CLKN_LVDS(0) => SP7_ZU_SPARE1N_CLKN_LVDS(0),
      SP7_ZU_SPARE1P_CLKP_LVDS(0) => SP7_ZU_SPARE1P_CLKP_LVDS(0),
      ZU_BOOT_STATUS_2V5 => ZU_BOOT_STATUS_2V5,
      ZU_DONE_2V5 => ZU_DONE_2V5,
      ZU_ERROR_OUT_2V5 => ZU_ERROR_OUT_2V5,
      ZU_ERROR_STATUS_2V5 => ZU_ERROR_STATUS_2V5,
      ZU_GNSS_1PPS => ZU_GNSS_1PPS,
      ZU_SP7_DMCU_RESET_STAT => ZU_SP7_DMCU_RESET_STAT,
      spi_rtl_0_io0_i => spi_rtl_0_io0_i,
      spi_rtl_0_io0_o => spi_rtl_0_io0_o,
      spi_rtl_0_io0_t => spi_rtl_0_io0_t,
      spi_rtl_0_io1_i => spi_rtl_0_io1_i,
      spi_rtl_0_io1_o => spi_rtl_0_io1_o,
      spi_rtl_0_io1_t => spi_rtl_0_io1_t,
      spi_rtl_0_io2_i => spi_rtl_0_io2_i,
      spi_rtl_0_io2_o => spi_rtl_0_io2_o,
      spi_rtl_0_io2_t => spi_rtl_0_io2_t,
      spi_rtl_0_io3_i => spi_rtl_0_io3_i,
      spi_rtl_0_io3_o => spi_rtl_0_io3_o,
      spi_rtl_0_io3_t => spi_rtl_0_io3_t,
      spi_rtl_0_ss_i(0) => spi_rtl_0_ss_i_0(0),
      spi_rtl_0_ss_o(0) => spi_rtl_0_ss_o_0(0),
      spi_rtl_0_ss_t => spi_rtl_0_ss_t
    );
spi_rtl_0_io0_iobuf: component IOBUF
     port map (
      I => spi_rtl_0_io0_o,
      IO => spi_rtl_0_io0_io,
      O => spi_rtl_0_io0_i,
      T => spi_rtl_0_io0_t
    );
spi_rtl_0_io1_iobuf: component IOBUF
     port map (
      I => spi_rtl_0_io1_o,
      IO => spi_rtl_0_io1_io,
      O => spi_rtl_0_io1_i,
      T => spi_rtl_0_io1_t
    );
spi_rtl_0_io2_iobuf: component IOBUF
     port map (
      I => spi_rtl_0_io2_o,
      IO => spi_rtl_0_io2_io,
      O => spi_rtl_0_io2_i,
      T => spi_rtl_0_io2_t
    );
spi_rtl_0_io3_iobuf: component IOBUF
     port map (
      I => spi_rtl_0_io3_o,
      IO => spi_rtl_0_io3_io,
      O => spi_rtl_0_io3_i,
      T => spi_rtl_0_io3_t
    );
spi_rtl_0_ss_iobuf_0: component IOBUF
     port map (
      I => spi_rtl_0_ss_o_0(0),
      IO => spi_rtl_0_ss_io(0),
      O => spi_rtl_0_ss_i_0(0),
      T => spi_rtl_0_ss_t
    );
end STRUCTURE;
